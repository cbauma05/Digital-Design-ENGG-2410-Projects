----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    13:38:00 10/31/2023 
-- Design Name: 
-- Module Name:    half_adder - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity half_adder is
    Port ( a_ha : in  STD_LOGIC;
           b_ha : in  STD_LOGIC;
           s_ha : out  STD_LOGIC;
           c_ha : out  STD_LOGIC);
end half_adder;

architecture Behavioral of half_adder is	
begin
	s_ha <= a_ha xor b_ha;
	c_ha <= a_ha and b_ha;

end Behavioral;

